//-------------------------------------------------------------------
//
//  COPYRIGHT (C) 2023, devin
//  balddonkey@outlook.com
//
//-------------------------------------------------------------------
//
//  Author      : Devin
//  Project		: project
//  Repository  : https://github.com/devindang/
//  Title       : file_name.v
//  Dependances : 
//  Editor      : VIM
//  Created     : 
//  Description : 
//
//-------------------------------------------------------------------

module file_name(

);


//------------------------ SIGNALS ------------------------//



//------------------------ PROCESS ------------------------//



//------------------------ INST ------------------------//


endmodule
