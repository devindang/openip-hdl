//-------------------------------------------------------------------
//
//  COPYRIGHT (C) 2023, devin
//  balddonkey@outlook.com
//
//-------------------------------------------------------------------
//
//  Author      : Devin
//  Project		: OPENIP-HDL
//  Repository  : https://github.com/devindang/openip-hdl
//  Title       : uart_clkdiv.v
//  Dependances : 
//  Editor      : VIM
//  Created     : 
//  Description : use PLL instead.
//
//-------------------------------------------------------------------

`include "uart_defines.v"

module uart_clkdiv(

);


//------------------------ SIGNALS ------------------------//



//------------------------ PROCESS ------------------------//



//------------------------ INST ------------------------//


endmodule